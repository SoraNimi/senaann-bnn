.PARAM mvdd=1.8
VVDD VDD 0 DC mvdd
VVREF VREF 0 DC mvdd
VVREFB VREFB 0 DC 0
vx0 x0 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx1 x1 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx2 x2 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx3 x3 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx4 x4 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx5 x5 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx6 x6 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx7 x7 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx8 x8 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx9 x9 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx10 x10 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx11 x11 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx12 x12 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx13 x13 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx14 x14 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx15 x15 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx16 x16 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx17 x17 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx18 x18 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx19 x19 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx20 x20 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx21 x21 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx22 x22 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx23 x23 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx24 x24 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx25 x25 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx26 x26 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx27 x27 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx28 x28 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx29 x29 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx30 x30 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx31 x31 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx32 x32 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx33 x33 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx34 x34 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx35 x35 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx36 x36 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx37 x37 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx38 x38 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx39 x39 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx40 x40 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx41 x41 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx42 x42 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx43 x43 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx44 x44 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx45 x45 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx46 x46 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx47 x47 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx48 x48 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx49 x49 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx50 x50 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx51 x51 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx52 x52 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx53 x53 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx54 x54 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx55 x55 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx56 x56 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx57 x57 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx58 x58 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx59 x59 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx60 x60 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx61 x61 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx62 x62 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx63 x63 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx64 x64 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx65 x65 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx66 x66 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx67 x67 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx68 x68 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx69 x69 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx70 x70 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx71 x71 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx72 x72 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx73 x73 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx74 x74 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx75 x75 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx76 x76 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx77 x77 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx78 x78 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx79 x79 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx80 x80 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx81 x81 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx82 x82 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx83 x83 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx84 x84 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx85 x85 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx86 x86 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx87 x87 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx88 x88 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx89 x89 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx90 x90 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx91 x91 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx92 x92 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx93 x93 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx94 x94 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx95 x95 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx96 x96 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx97 x97 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx98 x98 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx99 x99 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx100 x100 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx101 x101 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx102 x102 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx103 x103 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx104 x104 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx105 x105 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx106 x106 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx107 x107 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx108 x108 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx109 x109 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx110 x110 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx111 x111 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx112 x112 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx113 x113 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx114 x114 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx115 x115 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx116 x116 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx117 x117 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx118 x118 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx119 x119 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx120 x120 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx121 x121 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx122 x122 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx123 x123 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx124 x124 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx125 x125 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx126 x126 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx127 x127 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx128 x128 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx129 x129 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx130 x130 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx131 x131 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx132 x132 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx133 x133 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx134 x134 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx135 x135 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx136 x136 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx137 x137 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx138 x138 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx139 x139 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx140 x140 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx141 x141 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx142 x142 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx143 x143 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx144 x144 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx145 x145 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx146 x146 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx147 x147 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx148 x148 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx149 x149 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx150 x150 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx151 x151 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx152 x152 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx153 x153 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx154 x154 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx155 x155 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx156 x156 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx157 x157 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx158 x158 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx159 x159 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx160 x160 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx161 x161 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx162 x162 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx163 x163 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx164 x164 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx165 x165 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx166 x166 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx167 x167 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx168 x168 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx169 x169 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx170 x170 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx171 x171 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx172 x172 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx173 x173 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx174 x174 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx175 x175 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx176 x176 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx177 x177 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx178 x178 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx179 x179 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx180 x180 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx181 x181 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx182 x182 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx183 x183 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx184 x184 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx185 x185 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx186 x186 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx187 x187 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx188 x188 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx189 x189 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx190 x190 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx191 x191 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx192 x192 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx193 x193 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx194 x194 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx195 x195 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx196 x196 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx197 x197 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx198 x198 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx199 x199 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx200 x200 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx201 x201 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx202 x202 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx203 x203 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx204 x204 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx205 x205 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx206 x206 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx207 x207 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx208 x208 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx209 x209 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx210 x210 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx211 x211 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx212 x212 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx213 x213 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx214 x214 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx215 x215 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx216 x216 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx217 x217 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx218 x218 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx219 x219 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx220 x220 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx221 x221 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx222 x222 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx223 x223 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx224 x224 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx225 x225 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx226 x226 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx227 x227 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx228 x228 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx229 x229 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx230 x230 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx231 x231 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx232 x232 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx233 x233 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx234 x234 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx235 x235 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx236 x236 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx237 x237 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx238 x238 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx239 x239 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx240 x240 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx241 x241 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx242 x242 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx243 x243 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx244 x244 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx245 x245 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx246 x246 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx247 x247 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx248 x248 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx249 x249 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx250 x250 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx251 x251 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx252 x252 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx253 x253 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx254 x254 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx255 x255 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx256 x256 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx257 x257 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx258 x258 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx259 x259 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx260 x260 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx261 x261 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx262 x262 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx263 x263 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx264 x264 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx265 x265 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx266 x266 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx267 x267 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx268 x268 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx269 x269 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx270 x270 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx271 x271 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx272 x272 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx273 x273 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx274 x274 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx275 x275 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx276 x276 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx277 x277 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx278 x278 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx279 x279 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx280 x280 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx281 x281 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx282 x282 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx283 x283 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx284 x284 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx285 x285 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx286 x286 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx287 x287 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx288 x288 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx289 x289 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx290 x290 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx291 x291 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx292 x292 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx293 x293 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx294 x294 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx295 x295 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx296 x296 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx297 x297 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx298 x298 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx299 x299 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx300 x300 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx301 x301 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx302 x302 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx303 x303 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx304 x304 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx305 x305 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx306 x306 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx307 x307 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx308 x308 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx309 x309 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx310 x310 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx311 x311 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx312 x312 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx313 x313 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx314 x314 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx315 x315 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx316 x316 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx317 x317 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx318 x318 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx319 x319 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx320 x320 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx321 x321 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx322 x322 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx323 x323 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx324 x324 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx325 x325 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx326 x326 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx327 x327 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx328 x328 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx329 x329 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx330 x330 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx331 x331 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx332 x332 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx333 x333 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx334 x334 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx335 x335 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx336 x336 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx337 x337 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx338 x338 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx339 x339 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx340 x340 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx341 x341 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx342 x342 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx343 x343 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx344 x344 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx345 x345 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx346 x346 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx347 x347 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx348 x348 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx349 x349 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx350 x350 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx351 x351 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx352 x352 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx353 x353 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx354 x354 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx355 x355 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx356 x356 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx357 x357 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx358 x358 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx359 x359 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx360 x360 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx361 x361 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx362 x362 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx363 x363 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx364 x364 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx365 x365 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx366 x366 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx367 x367 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx368 x368 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx369 x369 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx370 x370 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx371 x371 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx372 x372 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx373 x373 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx374 x374 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx375 x375 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx376 x376 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx377 x377 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx378 x378 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx379 x379 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx380 x380 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx381 x381 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx382 x382 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx383 x383 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx384 x384 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx385 x385 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx386 x386 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx387 x387 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx388 x388 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx389 x389 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx390 x390 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx391 x391 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx392 x392 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx393 x393 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx394 x394 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx395 x395 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx396 x396 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx397 x397 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx398 x398 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx399 x399 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx400 x400 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx401 x401 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx402 x402 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx403 x403 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx404 x404 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx405 x405 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx406 x406 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx407 x407 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx408 x408 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx409 x409 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx410 x410 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx411 x411 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx412 x412 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx413 x413 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx414 x414 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx415 x415 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx416 x416 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx417 x417 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx418 x418 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx419 x419 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx420 x420 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx421 x421 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx422 x422 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx423 x423 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx424 x424 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx425 x425 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx426 x426 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx427 x427 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx428 x428 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx429 x429 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx430 x430 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx431 x431 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx432 x432 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx433 x433 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx434 x434 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx435 x435 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx436 x436 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx437 x437 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx438 x438 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx439 x439 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx440 x440 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx441 x441 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx442 x442 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx443 x443 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx444 x444 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx445 x445 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx446 x446 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx447 x447 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx448 x448 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx449 x449 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx450 x450 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx451 x451 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx452 x452 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx453 x453 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx454 x454 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx455 x455 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx456 x456 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx457 x457 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx458 x458 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx459 x459 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx460 x460 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx461 x461 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx462 x462 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx463 x463 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx464 x464 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx465 x465 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx466 x466 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx467 x467 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx468 x468 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx469 x469 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx470 x470 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx471 x471 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx472 x472 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx473 x473 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx474 x474 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx475 x475 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx476 x476 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx477 x477 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx478 x478 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx479 x479 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx480 x480 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx481 x481 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx482 x482 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx483 x483 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx484 x484 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx485 x485 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx486 x486 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx487 x487 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx488 x488 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx489 x489 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx490 x490 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx491 x491 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx492 x492 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx493 x493 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx494 x494 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx495 x495 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx496 x496 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx497 x497 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx498 x498 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx499 x499 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx500 x500 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx501 x501 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx502 x502 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx503 x503 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx504 x504 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx505 x505 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx506 x506 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx507 x507 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx508 x508 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx509 x509 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx510 x510 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx511 x511 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx512 x512 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx513 x513 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx514 x514 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx515 x515 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx516 x516 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx517 x517 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx518 x518 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx519 x519 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx520 x520 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx521 x521 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx522 x522 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx523 x523 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx524 x524 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx525 x525 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx526 x526 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx527 x527 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx528 x528 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx529 x529 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx530 x530 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx531 x531 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx532 x532 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx533 x533 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx534 x534 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx535 x535 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx536 x536 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx537 x537 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx538 x538 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx539 x539 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx540 x540 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx541 x541 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx542 x542 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx543 x543 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx544 x544 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx545 x545 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx546 x546 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx547 x547 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx548 x548 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx549 x549 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx550 x550 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx551 x551 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx552 x552 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx553 x553 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx554 x554 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx555 x555 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx556 x556 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx557 x557 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx558 x558 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx559 x559 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx560 x560 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx561 x561 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx562 x562 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx563 x563 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx564 x564 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx565 x565 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx566 x566 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx567 x567 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx568 x568 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx569 x569 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx570 x570 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx571 x571 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx572 x572 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx573 x573 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx574 x574 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx575 x575 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx576 x576 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx577 x577 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx578 x578 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx579 x579 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx580 x580 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx581 x581 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx582 x582 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx583 x583 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx584 x584 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx585 x585 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx586 x586 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx587 x587 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx588 x588 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx589 x589 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx590 x590 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx591 x591 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx592 x592 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx593 x593 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx594 x594 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx595 x595 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx596 x596 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx597 x597 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx598 x598 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx599 x599 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx600 x600 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx601 x601 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx602 x602 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx603 x603 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx604 x604 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx605 x605 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx606 x606 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx607 x607 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx608 x608 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx609 x609 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx610 x610 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx611 x611 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx612 x612 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx613 x613 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx614 x614 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx615 x615 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx616 x616 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx617 x617 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx618 x618 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx619 x619 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx620 x620 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx621 x621 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx622 x622 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx623 x623 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx624 x624 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx625 x625 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx626 x626 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx627 x627 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx628 x628 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx629 x629 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx630 x630 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx631 x631 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx632 x632 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx633 x633 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx634 x634 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx635 x635 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx636 x636 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx637 x637 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx638 x638 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx639 x639 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx640 x640 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx641 x641 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx642 x642 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx643 x643 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx644 x644 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx645 x645 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx646 x646 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx647 x647 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx648 x648 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx649 x649 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx650 x650 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx651 x651 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx652 x652 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx653 x653 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx654 x654 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx655 x655 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx656 x656 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx657 x657 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx658 x658 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx659 x659 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx660 x660 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx661 x661 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx662 x662 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx663 x663 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx664 x664 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx665 x665 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx666 x666 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx667 x667 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx668 x668 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx669 x669 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx670 x670 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx671 x671 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx672 x672 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx673 x673 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx674 x674 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx675 x675 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx676 x676 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx677 x677 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx678 x678 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx679 x679 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx680 x680 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx681 x681 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx682 x682 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx683 x683 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx684 x684 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx685 x685 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx686 x686 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx687 x687 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx688 x688 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx689 x689 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx690 x690 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx691 x691 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx692 x692 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx693 x693 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx694 x694 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx695 x695 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx696 x696 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx697 x697 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx698 x698 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx699 x699 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx700 x700 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx701 x701 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx702 x702 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx703 x703 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx704 x704 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx705 x705 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx706 x706 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx707 x707 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx708 x708 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx709 x709 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx710 x710 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx711 x711 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx712 x712 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx713 x713 0 PWL  
+	0n		mvdd
+	20n		mvdd
+	25n	    mvdd
+	200n    mvdd

vx714 x714 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx715 x715 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx716 x716 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx717 x717 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx718 x718 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx719 x719 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx720 x720 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx721 x721 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx722 x722 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx723 x723 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx724 x724 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx725 x725 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx726 x726 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx727 x727 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx728 x728 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx729 x729 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx730 x730 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx731 x731 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx732 x732 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx733 x733 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx734 x734 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx735 x735 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx736 x736 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx737 x737 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx738 x738 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx739 x739 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx740 x740 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx741 x741 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx742 x742 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx743 x743 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx744 x744 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx745 x745 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx746 x746 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx747 x747 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx748 x748 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx749 x749 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx750 x750 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx751 x751 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx752 x752 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx753 x753 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx754 x754 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx755 x755 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx756 x756 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx757 x757 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx758 x758 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx759 x759 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx760 x760 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx761 x761 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx762 x762 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx763 x763 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx764 x764 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx765 x765 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx766 x766 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx767 x767 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx768 x768 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx769 x769 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx770 x770 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx771 x771 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx772 x772 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx773 x773 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx774 x774 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx775 x775 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx776 x776 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx777 x777 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx778 x778 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx779 x779 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx780 x780 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx781 x781 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx782 x782 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

vx783 x783 0 PWL  
+	0n		0
+	20n		0
+	25n	    0
+	200n    0

.END
